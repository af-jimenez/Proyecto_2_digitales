LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE work.my_pkg.ALL;
----------------------------------------
ENTITY main_FSM IS
	PORT	(	clk				:	IN	STD_LOGIC;
				rst				:	IN	STD_LOGIC;
				ena				:	IN	STD_LOGIC;
				str_btn			:	IN	STD_LOGIC;
				col_izq			:	IN	STD_LOGIC;
				col_der			:	IN	STD_LOGIC;
				max_izq			:	IN	STD_LOGIC;
				max_der			:	IN	STD_LOGIC;
				tick_timer_1s	:	IN	STD_LOGIC;
				tick_timer_3s	:	IN	STD_LOGIC;
				tick_timer_g	:	IN	STD_LOGIC;
				tick_timer_w	:	IN	STD_LOGIC;
				timer_ena_3s	:	OUT	STD_LOGIC	:=	'0';
				timer_ena_g		:	OUT	STD_LOGIC	:=	'0';
				timer_ena_w		:	OUT	STD_LOGIC	:=	'0';
				goal_sig_1		:	OUT	STD_LOGIC	:=	'0';
				goal_sig_2		:	OUT	STD_LOGIC	:=	'0';
				rst_game			:	OUT	STD_LOGIC	:=	'1';
				wr_en				:	OUT	STD_LOGIC;
				w_addr_j			:	OUT	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
				w_addr_i			:	OUT	STD_LOGIC_VECTOR( 2 DOWNTO 0 );
				w_data			:	OUT	STD_LOGIC);
END ENTITY;
----------------------------------------
ARCHITECTURE arch OF main_FSM IS
	
	SIGNAL	w_addr_s0_j	:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
	SIGNAL	w_addr_s0_i	:	STD_LOGIC_VECTOR( 2 DOWNTO 0 );
	SIGNAL	w_data_s0	:	STD_LOGIC;
	SIGNAL	wr_en_s0		:	STD_LOGIC;
	SIGNAL	w_addr_s1_j	:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
	SIGNAL	w_addr_s1_i	:	STD_LOGIC_VECTOR( 2 DOWNTO 0 );
	SIGNAL	w_data_s1	:	STD_LOGIC;
	SIGNAL	wr_en_s1		:	STD_LOGIC;
	SIGNAL	w_addr_s3_j	:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
	SIGNAL	w_addr_s3_i	:	STD_LOGIC_VECTOR( 2 DOWNTO 0 );
	SIGNAL	w_data_s3	:	STD_LOGIC;
	SIGNAL	wr_en_s3		:	STD_LOGIC;
	SIGNAL	w_addr_s4_j	:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
	SIGNAL	w_addr_s4_i	:	STD_LOGIC_VECTOR( 2 DOWNTO 0 );
	SIGNAL	w_data_s4	:	STD_LOGIC;
	SIGNAL	wr_en_s4		:	STD_LOGIC;
	SIGNAL	w_addr_s6_j	:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
	SIGNAL	w_addr_s6_i	:	STD_LOGIC_VECTOR( 2 DOWNTO 0 );
	SIGNAL	w_data_s6	:	STD_LOGIC;
	SIGNAL	wr_en_s6		:	STD_LOGIC;
	SIGNAL	w_addr_sc_j	:	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
	SIGNAL	w_addr_sc_i	:	STD_LOGIC_VECTOR( 2 DOWNTO 0 );
	SIGNAL	w_data_sc	:	STD_LOGIC;
	SIGNAL	wr_en_sc		:	STD_LOGIC;
	
	SIGNAL	anim_imgs	:	imgs_mtx( 0 TO 3 );
	SIGNAL	anim_img	:	img_mtx;

	
	TYPE state IS (st0, st1, st2, st3, st4, st5, st6, st7);
	SIGNAL pr_state, nx_state	:	state;
	
BEGIN
	
	anim_imgs(0)	<= (	conv_slv("0000000000000000"),
							conv_slv("0111011101110111"),
							conv_slv("0001010101010101"),
							conv_slv("0111010101010101"),
							conv_slv("0101010101010111"),
							conv_slv("0101010101010001"),
							conv_slv("0111010101110001"),
							conv_slv("0000000000000000"));
	
	anim_imgs(1)	<= (	conv_slv("0000000000000000"),
							conv_slv("0001011101110111"),
							conv_slv("0001010101010001"),
							conv_slv("0001011101010111"),
							conv_slv("0001010101010101"),
							conv_slv("0001010101010101"),
							conv_slv("0111010101110111"),
							conv_slv("0000000000000000"));
	
	anim_imgs(2)	<= (	conv_slv("0000000000000000"),
							conv_slv("0001000000111100"),
							conv_slv("0001100000100100"),
							conv_slv("0001010000100100"),
							conv_slv("0001000000111100"),
							conv_slv("0001000000000100"),
							conv_slv("0011100000000100"),
							conv_slv("0000000000000000"));
	
	anim_imgs(3)	<= (	conv_slv("0000000000000000"),
							conv_slv("0011100000111100"),
							conv_slv("0010000000100100"),
							conv_slv("0011100000100100"),
							conv_slv("0000100000111100"),
							conv_slv("0000100000000100"),
							conv_slv("0011100000000100"),
							conv_slv("0000000000000000"));
	
	pong_print:	ENTITY work.imageManagement
				PORT MAP(clk      =>	clk,
						rst      =>	rst,
						ena      =>	ena,
						imageIn	=>	anim_imgs(0),
						wr_en		=>	wr_en_s0,
						w_addr_j	=>	w_addr_s0_j,
						w_addr_i	=>	w_addr_s0_i,
						w_data	=>	w_data_s0);
	
	conteo_fsm: ENTITY work.countdown_FSM
				PORT MAP(clk     		=>	clk,
						rst      		=>	rst,
						ena      		=>	ena,
						tick_timer_1s	=>	tick_timer_1s,
						wr_en			=>	wr_en_s1,
						w_addr_j		=>	w_addr_s1_j,
						w_addr_i		=>	w_addr_s1_i,
						w_data			=>	w_data_s1);
	
	g_print:	ENTITY work.imageManagement
				PORT MAP(clk      =>	clk,
						rst      =>	rst,
						ena      =>	ena,
						imageIn	=>	anim_imgs(1),
						wr_en		=>	wr_en_s3,
						w_addr_j	=>	w_addr_s3_j,
						w_addr_i	=>	w_addr_s3_i,
						w_data	=>	w_data_s3);
	
	w1_print:	ENTITY work.imageManagement
				PORT MAP(clk      =>	clk,
						rst      =>	rst,
						ena      =>	ena,
						imageIn	=>	anim_imgs(2),
						wr_en		=>	wr_en_s4,
						w_addr_j	=>	w_addr_s4_j,
						w_addr_i	=>	w_addr_s4_i,
						w_data	=>	w_data_s4);
	
	w2_print:	ENTITY work.imageManagement
				PORT MAP(clk      =>	clk,
						rst      =>	rst,
						ena      =>	ena,
						imageIn	=>	anim_imgs(3),
						wr_en		=>	wr_en_s6,
						w_addr_j	=>	w_addr_s6_j,
						w_addr_i	=>	w_addr_s6_i,
						w_data	=>	w_data_s6);
	
	anim_img		<= (	conv_slv("0000000000000000"),
							conv_slv("0000000000000000"),
							conv_slv("0000000000000000"),
							conv_slv("0000000000000000"),
							conv_slv("0000000000000000"),
							conv_slv("0000000000000000"),
							conv_slv("0000000000000000"),
							conv_slv("0000000000000000"));
	
	framec_print: ENTITY work.imageManagement
				PORT MAP (clk      =>	clk,
							rst      =>	rst,
							ena      =>	'1',
							imageIn	=>	anim_img,
							wr_en		=>	wr_en_sc,
							w_addr_j	=>	w_addr_sc_j,
							w_addr_i	=>	w_addr_sc_i,
							w_data	=>	w_data_sc);
	
	-------------------------------------------------------------
	--                 LOWER SECTION OF FSM                    --
	-------------------------------------------------------------
	sequential: PROCESS(rst, clk)
	BEGIN
		IF (rst = '1') THEN
			pr_state	<=	st0;
		ELSIF (rising_edge(clk)) THEN
			pr_state	<=	nx_state;
		END IF;
	END PROCESS sequential;
	
	-------------------------------------------------------------
	--                 UPPER SECTION OF FSM                    --
	-------------------------------------------------------------
	combinational: PROCESS(str_btn, col_der, col_izq, max_der, max_izq, tick_timer_3s, tick_timer_1s, tick_timer_g, tick_timer_w)
	BEGIN
		CASE pr_state IS
			WHEN st0	=>
				
				wr_en		<=	wr_en_s0;
				w_addr_j	<=	w_addr_s0_j;
				w_addr_i	<=	w_addr_s0_i;
				w_data	<=	w_data_s0;
					
				timer_ena_3s	<=	'0';
				timer_ena_g		<=	'0';
				timer_ena_w		<=	'0';
				rst_game		<=	'1';
				
				goal_sig_1	<=	'0';
				goal_sig_2	<=	'0';
				
				IF (str_btn = '1') THEN
					nx_state	<= st7;
				ELSE
					nx_state	<= st0;
				END IF;
			WHEN st1	=>
				
				timer_ena_3s	<=	'1';
				timer_ena_g		<=	'0';
				timer_ena_w		<=	'0';
				rst_game		<=	'1';
				
				wr_en		<=	wr_en_s1;
				w_addr_j	<=	w_addr_s1_j;
				w_addr_i	<=	w_addr_s1_i;
				w_data	<=	w_data_s1;
				
				goal_sig_1	<=	'0';
				goal_sig_2	<=	'0';
				
				IF (tick_timer_3s = '1') THEN
					nx_state	<= st2;
				ELSE
					nx_state	<= st1;
				END IF;
			WHEN st2	=>
				
				wr_en		<=	'1';
				w_addr_j	<=	"0000";
				w_addr_i	<=	"000";
				w_data	<=	'0';
				
				timer_ena_3s	<=	'0';
				timer_ena_g		<=	'0';
				timer_ena_w		<=	'0';
				rst_game		<=	'0';
				
				IF (col_der = '1') THEN
					nx_state	<= st3;	
				ELSIF (col_izq = '1') THEN
					nx_state	<= st5;
				ELSIF (max_der = '1') THEN
					nx_state	<= st4;
				ELSIF (max_izq = '1') THEN
					nx_state	<= st6;
				ELSE
					nx_state	<= st2;
				END IF;
				
			WHEN st3	=>
				
				wr_en		<=	wr_en_s3;
				w_addr_j	<=	w_addr_s3_j;
				w_addr_i	<=	w_addr_s3_i;
				w_data	<=	w_data_s3;
				
				timer_ena_3s	<=	'0';
				timer_ena_g		<=	'1';
				timer_ena_w		<=	'0';
				rst_game		<=	'1';
				
				goal_sig_1	<=	'1';
				goal_sig_2	<=	'0';
					
				IF (max_der = '1') THEN
					nx_state	<= st4;
				ELSIF (tick_timer_g = '1') THEN
					nx_state	<= st2;
				ELSE
					nx_state	<= st3;
				END IF;
				
			WHEN st4	=>
				
				wr_en		<=	wr_en_s4;
				w_addr_j	<=	w_addr_s4_j;
				w_addr_i	<=	w_addr_s4_i;
				w_data	<=	w_data_s4;
				
				timer_ena_3s	<=	'0';
				timer_ena_g		<=	'0';
				timer_ena_w		<=	'1';
				rst_game		<=	'1';
				
				goal_sig_1	<=	'0';
				goal_sig_2	<=	'0';
				
				IF (tick_timer_w = '1') THEN
					nx_state	<= st0;
				ELSE
					nx_state	<= st4;
				END IF;
				
			WHEN st5	=>
				
				wr_en		<=	wr_en_s3;
				w_addr_j	<=	w_addr_s3_j;
				w_addr_i	<=	w_addr_s3_i;
				w_data	<=	w_data_s3;
				
				timer_ena_3s	<=	'0';
				timer_ena_g		<=	'1';
				timer_ena_w		<=	'0';
				rst_game		<=	'1';
				
				IF (max_izq = '1') THEN
					nx_state	<= st6;
				ELSIF (tick_timer_g = '1') THEN
					nx_state	<= st2;
				ELSE
					nx_state	<= st5;
				END IF;
			
				goal_sig_2	<=	'1';
				goal_sig_1	<=	'0';
			
			WHEN st6	=>
				
				wr_en		<=	wr_en_s6;
				w_addr_j	<=	w_addr_s6_j;
				w_addr_i	<=	w_addr_s6_i;
				w_data	<=	w_data_s6;
					
				timer_ena_3s	<=	'0';
				timer_ena_g		<=	'0';
				timer_ena_w		<=	'1';
				rst_game		<=	'1';
				
				goal_sig_1	<=	'0';
				goal_sig_2	<=	'0';
					
				IF (tick_timer_w = '1') THEN
					nx_state	<= st0;
				ELSE
					nx_state	<= st6;
				END IF;
				WHEN st7	=>
				wr_en		<=	wr_en_sc;
				w_addr_j	<=	w_addr_sc_j;
				w_addr_i	<=	w_addr_sc_i;
				w_data	<=	w_data_sc;
				nx_state	<=	st1;
		END CASE;
	END PROCESS combinational;
END ARCHITECTURE;